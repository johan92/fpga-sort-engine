`ifndef _SORT_DEFINES_SVH__
`define _SORT_DEFINES_SVH__


typedef enum { 
               RANDOM,
               INCREASING,
               DECREASING,
               CONSTANT
             } sort_trans_type_t;

`endif // _SORT_DEFINES_SVH__

