package sort_tb;

// including in order
`include "sort_defines.svh"
`include "sort_trans.sv"
`include "sort_driver.sv"
`include "sort_generator.sv"
`include "sort_monitor.sv"
`include "sort_scoreboard.sv"
`include "sort_environment.sv"

endpackage
